.title KiCad schematic
.include "C:/AE/ZXCT1010/_models/BZX84C4V7.spice.txt"
.include "C:/AE/ZXCT1010/_models/C2012C0G2A102J060AA_p.mod"
.include "C:/AE/ZXCT1010/_models/CGJ4C2C0G2A101J060AA_p.mod"
.include "C:/AE/ZXCT1010/_models/FMMT597.spice.txt"
.include "C:/AE/ZXCT1010/_models/SMAZ15.spice.txt"
.include "C:/AE/ZXCT1010/_models/ZXCT1010.spice.txt"
V1 /PWR_IN 0 {VSOURCE}
R3 /BASE 0 {RBASE}
R1 /OUT /FILTER {RFILTER}
XU2 /OUT 0 C2012C0G2A102J060AA_p
Q1 /FILTER /BASE /COCM FMMT597
XU1 0 /OUT DI_BZX84C4V7
R2 /FILTER 0 {RSET1}
R4 /FILTER 0 {RSET2}
R7 /PWR_IN /PWR_OUT {RSENSE1}
R8 /PWR_IN /PWR_OUT {RSENSE2}
R6 /PWR_OUT /SN {RLIM}
XU3 /BASE /PWR_IN SMAZ15
XU4 0 /COCM /PWR_IN /SN ZXCT1010
I1 /PWR_OUT 0 {ILOAD}
XU5 /PWR_IN /SN CGJ4C2C0G2A101J060AA_p
.end
